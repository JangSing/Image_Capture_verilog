`timescale 1ps/1ps

module I2C_CCD_Config_tb();	
input			iCLK;
input			iRST_N;
input 			iZOOM_MODE_SW;
output		I2C_SCLK;
inout		I2C_SDAT;
input 		iEXPOSURE_ADJ;
input		iEXPOSURE_DEC_p;	



endmodule